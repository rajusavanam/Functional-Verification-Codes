typedef uvm_sequencer #(tx) sequencer;
