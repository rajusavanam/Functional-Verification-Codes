typedef uvm_sequencer#(rd_tx)async_fifo_rd_sqr;
