`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "mem_design.sv"
`include "mem_assert.sv"
`include "mem_common.sv"
`include "mem_intfc.sv"
`include "mem_tx.sv"
`include "mem_sqr.sv"
`include "mem_seq_lib.sv"
`include "mem_drv.sv"
`include "mem_mon.sv"
`include "mem_cov.sv"
`include "mem_agent.sv"
`include "mem_sbd.sv"
`include "mem_env.sv"
`include "test_lib.sv"
`include "top.sv"
