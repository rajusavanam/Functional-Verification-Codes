`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "async_fifo_common.sv"
`include "async_fifo_intfc.sv"
`include "async_fifo_gray.v"

`include "wr_tx.sv"
`include "wr_seq_lib.sv"
`include "async_fifo_wr_sqr.sv"
`include "async_fifo_wr_drv.sv"
`include "async_fifo_wr_mon.sv"
`include "async_fifo_wr_cov.sv"
`include "async_fifo_wr_agent.sv"

`include "rd_tx.sv"
`include "rd_seq_lib.sv"
`include "async_fifo_rd_sqr.sv"
`include "async_fifo_rd_drv.sv"
`include "async_fifo_rd_mon.sv"
`include "async_fifo_rd_cov.sv"
`include "async_fifo_rd_agent.sv"


`include "async_fifo_sbd.sv"
`include "top_sqr.sv"
`include "top_seq_lib.sv"
`include "async_fifo_env.sv"
`include "test_lib.sv"
`include "top.sv"