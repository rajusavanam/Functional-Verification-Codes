`include "sy_fifo_intfc.sv"
`include "sy_fifo_common.sv"
`include "sync_fifo_design.v"
`include "sy_fifo_tx.sv"
`include "sy_fifo_gen.sv"
`include "sy_fifo_bfm.sv"
`include "sy_fifo_agent.sv"
`include "sy_fifo_env.sv"
`include "top.sv"
