typedef uvm_sequencer #(wr_tx)async_fifo_wr_sqr;
