typedef uvm_sequencer#(mem_tx)mem_sqr;
// The above line is same as below code. As usual all the common phases will be automatically called.

//class mem_sqr extends uvm_sequencer#(mem_tx);
//	`uvm_component_utils(mem_sqr)
//	`NEW_COMP
//endclass
