`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "common.sv"
`include "tx.sv"
`include "sequencer.sv"
`include "seq_lib.sv"
`include "driver.sv"
`include "coverage.sv"
`include "monitor.sv"
`include "agent.sv"
`include "sbd.sv"
`include "env.sv"
`include "test_lib.sv"
`include "top.sv"
