`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "axi_common.sv"
`include "axi_intf.sv"
`include "axi_tx.sv"
`include "axi_seq_lib.sv"
`include "axi_sequencer.sv"
`include "axi_driver.sv"
`include "axi_monitor.sv"
//`include "axi_mon_inorder.sv"
`include "axi_coverage.sv"
`include "axi_responder.sv"
`include "axi_agent.sv"
`include "axi_sbd.sv"
`include "axi_env.sv"
`include "axi_test_lib.sv"
`include "top.sv"
